library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

PACKAGE MY IS
	PROCEDURE square(
		SIGNAL Xcur,Ycur,Xpos,Ypos	:	IN INTEGER;
		SIGNAL RGB						:	OUT STD_LOGIC_VECTOR(3 downto 0);  --not much better color resolution with 8 bits hence 4 bits
		SIGNAL DRAW						: 	OUT STD_LOGIC
	);
END MY;

PACKAGE BODY MY IS
	PROCEDURE square(
		SIGNAL Xcur,Ycur,Xpos,Ypos:IN INTEGER;
		SIGNAL RGB:OUT STD_LOGIC_VECTOR(3 downto 0);
		SIGNAL DRAW: OUT STD_LOGIC) IS
	BEGIN
		IF(Xcur>Xpos AND Xcur<(Xpos+100) AND Ycur>Ypos AND Ycur<(Ypos+100))THEN
			RGB <= "1111";
			DRAW <= '1';
		ELSE
			DRAW <= '0';
		END IF;
	 
	END square;
END MY;